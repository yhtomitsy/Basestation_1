#include <orcapp_head>

module USERNAME_sig_delay (
  input wire   clk,
  input wire   rstn,
  input wire   in, 
  output wire  out
);

endmodule
