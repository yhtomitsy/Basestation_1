#include <orcapp_head>

module USERNAME_tinit_count (
  input wire    clk	,
  input wire    resetn	,
  output wire   tinit_done_o
);

endmodule

