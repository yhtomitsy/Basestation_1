#include <orcapp_head>

module USERNAME_dphy_2_cmos_ip #(
    parameter RX_TYPE      = "DSI",        // "DSI" or "CSI2" 
    parameter TX_TYPE      = "CMOS",       // "DSI", "CSI2", "CMOS" or "LVDS"
    parameter NUM_RX_LANE  = 4,            // 1, 2, 3 or 4
    parameter RX_GEAR      = 16,           // 8 or 16
    parameter DPHY_RX_IP   = "MIXEL",      // "MIXEL" or "LATTICE"
    parameter DATA_TYPE    = "RGB888",     // "RGB666", "RGB666_LOOSE", "RGB888", "RAW8", "RAW10", "RAW12", "YUV420-8", "LEGACY_YUV420_8",
                                           // "YUV420_8_CSPS", "YUV422_8", "YUV420_10", "YUV420_10_CSPS", "YUV420_10_CSPS" or "YUV422_10"
    parameter NUM_TX_CH    = 1,            // 1 or 2
    parameter PD_BUS_WIDTH = 24,           // 8, 10, 12, 18, 24, 36 or 48
    parameter RX_CLK_MODE  = "HS_LP",      // "HS_LP" or "HS_ONLY"
    parameter TX_WAIT_TIME = "LESS_15MS",  // "OVER_15MS" or "LESS_15MS"
    parameter LANE_ALIGN   = "OFF",         // Enable/Disable lane aligner
    parameter BYTECLK_MHZ  = 111,          // Target byte clock frequency
    parameter FIFO_DEPTH   = 16,           // Lane aligner FIFO depth
    parameter FIFO_TYPE0   = "EBR",        // Lane aligner FIFO type for lane 0
    parameter FIFO_TYPE1   = "EBR",        // Lane aligner FIFO type for lane 1
    parameter FIFO_TYPE2   = "EBR",        // Lane aligner FIFO type for lane 2
    parameter FIFO_TYPE3   = "EBR"         // Lane aligner FIFO type for lane 3
)
(
    input  wire                              reset_n_i,         // Reset, active low
    input  wire                              reset_lp_n_i,      // Reset to FFs using clk_lp_ctrl_i, active low
    input  wire                              reset_byte_n_i,    // Reset to FFs using clk_byte, active low
    input  wire                              reset_byte_fr_n_i, // Reset to FFs using clk_byte_fr_i, active low
    input  wire                              reset_pixel_n_i,   // Reset to FFs using clk_pixel_i, active low
    input  wire                              clk_lp_ctrl_i,     // clock to LP HS Controller on CLK lane
    input  wire                              clk_byte_fr_i,     // continuous byte clock, could be clk_byte_o/clk_byte_hs/refclk
    input  wire                              clk_pixel_i,       // pixel clock from PLL
    input  wire                              pll_lock_i,        // PLL lock indicator, active high; set to 1 if PLL is not in use

    ///// MIPI I/F
    inout  wire                              clk_p_i,           // DPHY clock (p)
    inout  wire                              clk_n_i,           // DPHY clock (n)
    inout  wire                              d0_p_io,           // DPHY D0 (p) in DSI
    inout  wire                              d0_n_io,           // DPHY D0 (n) in DSI
#ifdef PP_NUM_RX_LANE_4
    inout  wire                              d0_p_i,            // DPHY D0 (p) in CSI-2
    inout  wire                              d0_n_i,            // DPHY D0 (n) in CSI-2
    inout  wire                              d1_p_i,            // DPHY D1 (p)
    inout  wire                              d1_n_i,            // DPHY D1 (n)
    inout  wire                              d2_p_i,            // DPHY D2 (p)
    inout  wire                              d2_n_i,            // DPHY D2 (n)
    inout  wire                              d3_p_i,            // DPHY D3 (p)
    inout  wire                              d3_n_i,            // DPHY D3 (n)
#endif
#ifdef PP_NUM_RX_LANE_2
    inout  wire                              d0_p_i,            // DPHY D0 (p) in CSI-2
    inout  wire                              d0_n_i,            // DPHY D0 (n) in CSI-2
    inout  wire                              d1_p_i,            // DPHY D1 (p)
    inout  wire                              d1_n_i,            // DPHY D1 (n)
#endif
#ifdef PP_NUM_RX_LANE_1
    inout  wire                              d0_p_i,            // DPHY D0 (p) in CSI-2
    inout  wire                              d0_n_i,            // DPHY D0 (n) in CSI-2
#endif
    output wire                              clk_byte_o,        // non-continuous byte clock
    output wire                              clk_byte_fr_o,     // continuous byte clock in HS_ONLY mode 

    ///// DSI Rx only I/F                                   
    output wire                              lp_d0_rx_p_o,      // LP Rx Data on D0 (p)
    output wire                              lp_d0_rx_n_o,      // LP Rx Data on D0 (n)
    output wire                              lp_d1_rx_p_o,      // LP Rx Data on D1 (p)
    output wire                              lp_d1_rx_n_o,      // LP Rx Data on D1 (n)
    output wire                              lp_d2_rx_p_o,      // LP Rx Data on D2 (p)
    output wire                              lp_d2_rx_n_o,      // LP Rx Data on D2 (n)
    output wire                              lp_d3_rx_p_o,      // LP Rx Data on D3 (p)
    output wire                              lp_d3_rx_n_o,      // LP Rx Data on D3 (n)
    output wire                              cd_d0_o,           // Contenion Detection on D0
    input  wire                              lp_d0_tx_en_i,     // LP Tx Data Enable on D0, active high
    input  wire                              lp_d0_tx_p_i,      // LP Tx Data on D0 (p)
    input  wire                              lp_d0_tx_n_i,      // LP Tx Data on D0 (n)

    ///// DSI to DSI only I/F
    output wire [RX_GEAR-1:0]                bd0_o,             // DPHY Byte Data 0
    output wire [RX_GEAR-1:0]                bd1_o,             // DPHY Byte Data 1
    output wire [RX_GEAR-1:0]                bd2_o,             // DPHY Byte Data 2
    output wire [RX_GEAR-1:0]                bd3_o,             // DPHY Byte Data 3

    ///// CSI-2 to CSI-2 only I/F (or potential customer use and/or debug signals)
    output wire                              sp_en_o,           // Short Packet Enable, active high
    output wire                              lp_en_o,           // Long Packet Enable, active high
    output wire [5:0]                        dt_o,              // Data Type    
    output wire [1:0]                        vc_o,              // Virtual Channel
    output wire [15:0]                       wc_o,              // Byte count
    output wire [NUM_RX_LANE*8-1:0]          bd_o,              // DPHY Byte Data (Gear8 only)

    ///// DSI to CMOS/FPD-LINK only I/F
    output wire                              vsync_o,           // Vertical Sync, active high
    output wire                              hsync_o,           // Horizontal Sync, active high
    output wire                              de_o,              // Data Enable, active high

    ///// DSI to FPD-LINK only I/F
    output wire [1:0]                        p_odd_o,           // Odd pixel indicator

    ///// CSI2 to CMOS only I/F
    output wire                              fv_o,              // Frame Valid, active high
    output wire                              lv_o,              // Line Valid, active high
 
    ///// CMOS/FPD-LINK Tx only I/F
//  output wire                              clk_pixel_o,       // Pixel Clock (center aligned)
    output wire [PD_BUS_WIDTH*NUM_TX_CH-1:0] pd_o,              // Pixel Data
    
    ///// Debug only outputs (or potential customer use)
    output wire                              term_clk_en_o,     // Termination Enable on CLK, active high
    output wire                              hs_d_en_o,         // HS mode Enable on D0, active high
    output wire [1:0]                        lp_hs_state_clk_o, // LP HS Controller (CLK) state machine
    output wire [1:0]                        lp_hs_state_d_o,   // LP HS Controller (D0) state machine
    output wire                              hs_sync_o,         // HS Sync, active high
    output wire                              capture_en_o,      // Capture Enable, active high
    output wire                              sp2_en_o,          // Short Packet Enable #2, active high
    output wire                              lp2_en_o,          // Long Packet Enable #2, active high
    output wire                              lp_av_en_o,        // Active Video Long Packet Enable, active high
    output wire                              lp2_av_en_o,       // Active Video Long Packet Enable #2, active high
    output wire [5:0]                        dt2_o,             // Data Type #2   
    output wire [1:0]                        vc2_o,             // Virtual Channel #2
    output wire [15:0]                       wc2_o,             // Byte count #2
    output wire [7:0]                        ecc_o,             // ECC of Packet Header #2   
    output wire [7:0]                        ecc2_o,            // ECC of Packet Header #2   
    output wire                              payload_en_o,      // Payload Enable, active high
    output wire [3:0]                        write_cycle_o,     // Payload Data Write Cycle
    output wire                              mem_we_o,          // Payload Data Write Enable, active high
    output wire                              mem_re_o,          // Payload Data Read Enable, active high
    output wire [1:0]                        read_cycle_o,      // Pixel Data Read Cycle
    output wire [2:0]                        mem_radr_o         // Pixel Data Read Address
);


///// Internal Parameter Setting /////

localparam DT = ((RX_TYPE == "DSI") && (DATA_TYPE == "RGB666")) ?           6'h1E :
                ((RX_TYPE == "DSI") && (DATA_TYPE == "RGB666_LOOSE")) ?     6'h2E :
                ((RX_TYPE == "DSI") && (DATA_TYPE == "RGB888")) ?           6'h3E :
                ((RX_TYPE == "CSI2") && (DATA_TYPE == "RGB888")) ?          6'h24 :
                ((RX_TYPE == "CSI2") && (DATA_TYPE == "RAW10")) ?           6'h2B :
                ((RX_TYPE == "CSI2") && (DATA_TYPE == "RAW12")) ?           6'h2C :
                ((RX_TYPE == "CSI2") && (DATA_TYPE == "RAW8")) ?            6'h2A :
                ((RX_TYPE == "CSI2") && (DATA_TYPE == "YUV420_8")) ?        6'h18 :
                ((RX_TYPE == "CSI2") && (DATA_TYPE == "LEGACY_YUV420_8")) ? 6'h1A :
                ((RX_TYPE == "CSI2") && (DATA_TYPE == "YUV420_8_CSPS")) ?   6'h1C :
                ((RX_TYPE == "CSI2") && (DATA_TYPE == "YUV422_8")) ?        6'h1E :
                ((RX_TYPE == "CSI2") && (DATA_TYPE == "YUV420_10")) ?       6'h19 :
                ((RX_TYPE == "CSI2") && (DATA_TYPE == "YUV420_10_CSPS")) ?  6'h1D :
                ((RX_TYPE == "CSI2") && (DATA_TYPE == "YUV422_10")) ?       6'h1F : 6'h3E;

// No need to use rx fifo since data is already transferred to free-running byte clok
// inside dphy_rx_wrap using multicycle registers
localparam RX_FIFO = "OFF";

wire                           clk_byte_hs;
wire                           term_d0_en_w, term_d1_en_w, term_d2_en_w, term_d3_en_w;
wire                           term_d1_en_temp_w, term_d2_en_temp_w, term_d3_en_temp_w;
wire                           hs_d1_en_w, hs_d2_en_w, hs_d3_en_w;
wire                           hs_d1_en_temp_w, hs_d2_en_temp_w, hs_d3_en_temp_w;
wire                           capture_en_pre;
wire [RX_GEAR-1:0]             bd0, bd1, bd2, bd3, bd0_pre, bd1_pre, bd2_pre, bd3_pre;
wire                           lp_clk_rx_p, lp_clk_rx_n;
wire                           lp_av_en, lp2_av_en;
wire [NUM_RX_LANE*RX_GEAR-1:0] payload;

// Encountered synthesis error when driving unused dphy lanes with 1
// net \dphy_2_cmos/pwr is constantly driven from multiple places at instance \dphy_2_cmos/dsi.dsi_rx/d_sot_det_3__I_0_33, on port DN2. VDB-1000
// Done: error code 2
//wire                           d1_p, d1_n, d2_p, d2_n, d3_p, d3_n;
//generate
//    assign  d1_p = (NUM_RX_LANE > 1) ? d1_p_i : 1'b1; 
//    assign  d1_n = (NUM_RX_LANE > 1) ? d1_n_i : 1'b1; 
//    assign  d2_p = (NUM_RX_LANE > 2) ? d2_p_i : 1'b1; 
//    assign  d2_n = (NUM_RX_LANE > 2) ? d2_n_i : 1'b1; 
//    assign  d3_p = (NUM_RX_LANE > 3) ? d3_p_i : 1'b1; 
//    assign  d3_n = (NUM_RX_LANE > 3) ? d3_n_i : 1'b1; 
//endgenerate

generate
    assign clk_byte_fr_o = (RX_CLK_MODE == "HS_ONLY") ? clk_byte_hs : 1'b0;
endgenerate

assign capture_en_o = capture_en_pre;
assign bd0_o = bd0_pre;
assign bd1_o = bd1_pre;
assign bd2_o = bd2_pre;
assign bd3_o = bd3_pre;

generate
    if (RX_TYPE == "DSI")
    begin : dsi
        USERNAME_dphy_rx_wrap
        dsi_rx (
            .reset_n_i        (reset_n_i),
            .reset_byte_n_i   (reset_byte_n_i),
            .reset_byte_fr_n_i(reset_byte_fr_n_i),
            .clk_byte_fr_i    (clk_byte_fr_i),
            .clk_p_i          (clk_p_i),
            .clk_n_i          (clk_n_i),
#ifdef PP_NUM_RX_LANE_4
            .d0_p_io          (d0_p_io),
            .d0_n_io          (d0_n_io),
            .d1_p_i           (d1_p_i),
            .d1_n_i           (d1_n_i),
            .d2_p_i           (d2_p_i),
            .d2_n_i           (d2_n_i),
            .d3_p_i           (d3_p_i),
            .d3_n_i           (d3_n_i),
#endif
#ifdef PP_NUM_RX_LANE_2
            .d0_p_io          (d0_p_io),
            .d0_n_io          (d0_n_io),
            .d1_p_i           (d1_p_i),
            .d1_n_i           (d1_n_i),
#endif
#ifdef PP_NUM_RX_LANE_1
            .d0_p_io          (d0_p_io),
            .d0_n_io          (d0_n_io),
#endif
            .term_clk_en_i    (term_clk_en_o),
            .term_d0_en_i     (term_d0_en_w),
            .term_d1_en_i     (term_d1_en_w),
            .term_d2_en_i     (term_d2_en_w),
            .term_d3_en_i     (term_d3_en_w),
            .hs_d0_en_i       (hs_d_en_o),
            .hs_d1_en_i       (hs_d1_en_w),
            .hs_d2_en_i       (hs_d2_en_w),
            .hs_d3_en_i       (hs_d3_en_w),
            .lp_d0_tx_en_i    (lp_d0_tx_en_i),
            .lp_d0_tx_p_i     (lp_d0_tx_p_i),
            .lp_d0_tx_n_i     (lp_d0_tx_n_i),

            .clk_hs_o         (clk_byte_hs), // byte clk output. used to clock hs_ctrl_d0
            .clk_byte_o       (clk_byte_o),  // used to latch data
            .bd0_o            (bd0),
            .bd1_o            (bd1),
            .bd2_o            (bd2),
            .bd3_o            (bd3),
            .hs_sync_o        (hs_sync_o),

            .lp_clk_rx_p_o    (lp_clk_rx_p),
            .lp_clk_rx_n_o    (lp_clk_rx_n),
            .lp_d0_rx_p_o     (lp_d0_rx_p_o),
            .lp_d0_rx_n_o     (lp_d0_rx_n_o),
            .lp_d1_rx_p_o     (lp_d1_rx_p_o),
            .lp_d1_rx_n_o     (lp_d1_rx_n_o),
            .lp_d2_rx_p_o     (lp_d2_rx_p_o),
            .lp_d2_rx_n_o     (lp_d2_rx_n_o),
            .lp_d3_rx_p_o     (lp_d3_rx_p_o),
            .lp_d3_rx_n_o     (lp_d3_rx_n_o),
            .cd_clk_o         (),
            .cd_d0_o          (cd_d0_o)
        );
    end
    else if (RX_TYPE == "CSI2")
    begin : csi2
        USERNAME_dphy_rx_wrap 
        csi_rx (
            .reset_n_i        (reset_n_i),
            .reset_byte_n_i   (reset_byte_n_i),
            .reset_byte_fr_n_i(reset_byte_fr_n_i),
            .clk_byte_fr_i    (clk_byte_fr_i),
            .clk_p_i          (clk_p_i),
            .clk_n_i          (clk_n_i),
#ifdef PP_NUM_RX_LANE_4
            .d0_p_io          (d0_p_i),
            .d0_n_io          (d0_n_i),
            .d1_p_i           (d1_p_i),
            .d1_n_i           (d1_n_i),
            .d2_p_i           (d2_p_i),
            .d2_n_i           (d2_n_i),
            .d3_p_i           (d3_p_i),
            .d3_n_i           (d3_n_i),
#endif
#ifdef PP_NUM_RX_LANE_2
            .d0_p_io          (d0_p_i),
            .d0_n_io          (d0_n_i),
            .d1_p_i           (d1_p_i),
            .d1_n_i           (d1_n_i),
#endif
#ifdef PP_NUM_RX_LANE_1
            .d0_p_io          (d0_p_i),
            .d0_n_io          (d0_n_i),
#endif
            .term_clk_en_i    (term_clk_en_o),
            .term_d0_en_i     (term_d0_en_w),
            .term_d1_en_i     (term_d1_en_w),
            .term_d2_en_i     (term_d2_en_w),
            .term_d3_en_i     (term_d3_en_w),
            .hs_d0_en_i       (hs_d_en_o),
            .hs_d1_en_i       (hs_d1_en_w),
            .hs_d2_en_i       (hs_d2_en_w),
            .hs_d3_en_i       (hs_d3_en_w),
            .lp_d0_tx_en_i    (1'b0),
            .lp_d0_tx_p_i     (1'b0),
            .lp_d0_tx_n_i     (1'b0),

            .clk_hs_o         (clk_byte_hs),
            .clk_byte_o       (clk_byte_o),
            .bd0_o            (bd0),
            .bd1_o            (bd1),
            .bd2_o            (bd2),
            .bd3_o            (bd3),
            .hs_sync_o        (hs_sync_o),

            .lp_clk_rx_p_o    (lp_clk_rx_p),
            .lp_clk_rx_n_o    (lp_clk_rx_n),
            .lp_d0_rx_p_o     (lp_d0_rx_p_o),
            .lp_d0_rx_n_o     (lp_d0_rx_n_o),
            .lp_d1_rx_p_o     (lp_d1_rx_p_o),
            .lp_d1_rx_n_o     (lp_d1_rx_n_o),
            .lp_d2_rx_p_o     (lp_d2_rx_p_o),
            .lp_d2_rx_n_o     (lp_d2_rx_n_o),
            .lp_d3_rx_p_o     (lp_d3_rx_p_o),
            .lp_d3_rx_n_o     (lp_d3_rx_n_o),
            .cd_clk_o         (),
            .cd_d0_o          (cd_d0_o)
        );
    end
endgenerate


USERNAME_rx_global_ctrl 
rx_global_ctrl (
    .reset_n_i         (reset_n_i),
    .reset_lp_n_i      (reset_lp_n_i),
    .reset_byte_fr_n_i (reset_byte_fr_n_i),
    .clk_lp_ctrl_i     (clk_lp_ctrl_i),
    .clk_byte_i        (clk_byte_o),
    .clk_byte_hs_i     (clk_byte_hs),
    .clk_byte_fr_i     (clk_byte_fr_i),// use stoppable byteclk clk_hs (clk_byte_fr_i),
    .pll_lock_i        (pll_lock_i),
    .bd0_i             (bd0),
    .bd1_i             (bd1),
    .bd2_i             (bd2),
    .bd3_i             (bd3),
    .lp_clk_p_i        (lp_clk_rx_p),
    .lp_clk_n_i        (lp_clk_rx_n),
    .lp_d0_p_i         (lp_d0_rx_p_o),
    .lp_d0_n_i         (lp_d0_rx_n_o),
    .lp_d1_p_i         (lp_d1_rx_p_o),
    .lp_d1_n_i         (lp_d1_rx_n_o),
    .lp_d2_p_i         (lp_d2_rx_p_o),
    .lp_d2_n_i         (lp_d2_rx_n_o),
    .lp_d3_p_i         (lp_d3_rx_p_o),
    .lp_d3_n_i         (lp_d3_rx_n_o),
    .hs_sync_i         (hs_sync_o),
    .bd0_o             (bd0_pre),
    .bd1_o             (bd1_pre),
    .bd2_o             (bd2_pre),
    .bd3_o             (bd3_pre),
    .term_clk_en_o     (term_clk_en_o),
    .term_d0_en_o      (term_d0_en_w),
    .hs_d0_en_o        (hs_d_en_o),
    .term_d1_en_o      (term_d1_en_temp_w),
    .hs_d1_en_o        (hs_d1_en_temp_w),
    .term_d2_en_o      (term_d2_en_temp_w),
    .hs_d2_en_o        (hs_d2_en_temp_w),
    .term_d3_en_o      (term_d3_en_temp_w),
    .hs_d3_en_o        (hs_d3_en_temp_w),
    .hs_sync_o         (capture_en_pre),
    .lp_hs_state_clk_o (lp_hs_state_clk_o),
    .lp_hs_state_d_o   (lp_hs_state_d_o)
);

// Workaround since LP data of lane 1,2,3 from Mixel is not correct
// Still checking if this is a Mixel bug or not
generate 
if (DPHY_RX_IP == "MIXEL") begin
  assign term_d1_en_w = term_d0_en_w;
  assign term_d2_en_w = term_d0_en_w;
  assign term_d3_en_w = term_d0_en_w;
  assign hs_d1_en_w   = hs_d_en_o;
  assign hs_d2_en_w   = hs_d_en_o;
  assign hs_d3_en_w   = hs_d_en_o;
end
else begin
  assign term_d1_en_w = term_d1_en_temp_w;
  assign term_d2_en_w = term_d2_en_temp_w;
  assign term_d3_en_w = term_d3_en_temp_w;
  assign hs_d1_en_w   = hs_d1_en_temp_w;
  assign hs_d2_en_w   = hs_d2_en_temp_w;
  assign hs_d3_en_w   = hs_d3_en_temp_w;
end
endgenerate

generate
    if ((RX_TYPE != "DSI") || (TX_TYPE != "DSI"))
    begin : non_DSI2DSI
        USERNAME_capture_ctrl 
        capture_ctrl (
            .reset_n_i      (reset_byte_fr_n_i),
            .clk_byte_i     (clk_byte_fr_i),
            .bd0_i          (bd0_pre),
            .bd1_i          (bd1_pre),
            .bd2_i          (bd2_pre),
            .bd3_i          (bd3_pre),
            .capture_en_i   (capture_en_pre),
            .sp_en_o        (sp_en_o),
            .sp2_en_o       (sp2_en_o),
            .lp_en_o        (lp_en_o),
            .lp_av_en_o     (lp_av_en_o),
            .lp2_en_o       (lp2_en_o),
            .lp2_av_en_o    (lp2_av_en_o),
            .payload_en_o   (payload_en_o),
            .payload_o      (payload),
            .bd_o           (bd_o),
            .vc_o           (vc_o),
            .vc2_o          (vc2_o),
            .wc_o           (wc_o),
            .wc2_o          (wc2_o),
            .dt_o           (dt_o),
            .dt2_o          (dt2_o),
            .ecc_o          (ecc_o),
            .ecc2_o         (ecc2_o)
        );
    end
endgenerate

generate
    if ((TX_TYPE == "CMOS") || (TX_TYPE == "LVDS"))
    begin : non_DPHY2DPHY
        USERNAME_byte2pixel 
        byte2pixel (
            .reset_byte_n_i  (reset_byte_fr_n_i),
            .reset_pixel_n_i (reset_pixel_n_i),
            .clk_byte_i      (clk_byte_fr_i),
            .clk_pixel_i     (clk_pixel_i),
            .sp_en_i         (sp_en_o),
            .sp2_en_i        (sp2_en_o),
            .dt_i            (dt_o),
            .dt2_i           (dt2_o),
            .lp_av_en_i      (lp_av_en_o),
            .lp2_av_en_i     (lp2_av_en_o),
            .payload_en_i    (payload_en_o),
            .payload_i       (payload),
            .wc_i            (wc_o),
            .wc2_i           (wc2_o),
            .vsync_o         (vsync_o),
            .hsync_o         (hsync_o),
            .fv_o            (fv_o),
            .lv_o            (lv_o),
            .de_o            (de_o),
            .pd_o            (pd_o),
            .p_odd_o         (p_odd_o),
            .write_cycle_o   (write_cycle_o),
            .mem_we_o        (mem_we_o),
            .mem_re_o        (mem_re_o),
            .read_cycle_o    (read_cycle_o),
            .mem_radr_o      (mem_radr_o)
        );
    end
endgenerate


endmodule
      
      
      
