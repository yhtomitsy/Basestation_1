`timescale 1 ns/1ps

module tracker_top_tb.v

end module

